package stimulus_pkg;

import uvm_pkg::*;

`include "env/packet.sv"
`include "env/packet_sequence.sv"

endpackage
