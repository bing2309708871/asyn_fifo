package test_pkg;

import uvm_pkg::*;
import stimulus_pkg::*;
import env_pkg::*;

`include "test/test_collection.sv"

endpackage
